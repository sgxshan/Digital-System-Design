library verilog;
use verilog.vl_types.all;
entity rxd_parity_vlg_vec_tst is
end rxd_parity_vlg_vec_tst;
