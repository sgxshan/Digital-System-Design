library verilog;
use verilog.vl_types.all;
entity rxd_shift_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        load            : in     vl_logic;
        reset           : in     vl_logic;
        rshift          : in     vl_logic;
        serial_in       : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end rxd_shift_vlg_sample_tst;
