library verilog;
use verilog.vl_types.all;
entity rxd_controller_vlg_vec_tst is
end rxd_controller_vlg_vec_tst;
