library verilog;
use verilog.vl_types.all;
entity rxd_shift_vlg_vec_tst is
end rxd_shift_vlg_vec_tst;
