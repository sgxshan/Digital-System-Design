library verilog;
use verilog.vl_types.all;
entity Inverter_vlg_vec_tst is
end Inverter_vlg_vec_tst;
