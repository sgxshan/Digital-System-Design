library verilog;
use verilog.vl_types.all;
entity Inverter_vlg_check_tst is
    port(
        txd             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Inverter_vlg_check_tst;
