library verilog;
use verilog.vl_types.all;
entity receiver_vlg_vec_tst is
end receiver_vlg_vec_tst;
