library verilog;
use verilog.vl_types.all;
entity IRtransceiver_vlg_vec_tst is
end IRtransceiver_vlg_vec_tst;
