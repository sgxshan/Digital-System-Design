library verilog;
use verilog.vl_types.all;
entity transmitter_vlg_vec_tst is
end transmitter_vlg_vec_tst;
