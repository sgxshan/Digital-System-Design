library verilog;
use verilog.vl_types.all;
entity baud_done_vlg_vec_tst is
end baud_done_vlg_vec_tst;
